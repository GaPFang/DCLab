module Block_Movement2Motor(
    
);

endmodule